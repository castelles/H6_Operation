library ieee;
use ieee.std_logic_1164.all;

entity div_freq is
	port (
			clk_50MHz  : in std_logic;	
			clk_1KHz	  : out std_logic
	);
end div_freq;

architecture arch of div_freq is
begin
	
end arch;