library ieee;
use ieee.std_logic_1164.all;

entity dsf_timer is
	port (
			clk       : in std_logic;
			trig   	 : in BIT;
			buz   	 : out BIT
	);
end dsf_timer;

architecture arch of dsf_timer is
begin
	
end arch;